*1BIT ADDER SUBCIRCUIT
.subckt 1bitadr 1 2 7 11 12 13
.include nand.cir
X1 1 2 3 13 nand
X2 1 3 4 13 nand
X3 3 2 5 13 nand
X4 4 5 6 13 nand
X5 6 7 8 13 nand
X6 6 8 9 13 nand
X7 8 7 10 13 nand
X8 9 10 11 13 nand
X9 8 3 12 13 nand
.ends 1bitadr
