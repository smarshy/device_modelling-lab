*1 BIT ADDER
.include nand.cir
X1 1 2 3 13 nand
X2 1 3 4 13 nand
X3 3 2 5 13 nand
X4 4 5 6 13 nand
X5 6 7 8 13 nand
X6 6 8 9 13 nand
X7 8 7 10 13 nand
X8 9 10 11 13 nand
X9 8 3 12 13 nand
Vdd 13 0 DC 5V
Va 1 0 PULSE (0 5 10n 0n 0n 25n 70n)
Vb 2 0 PULSE (0 5 5n 0n 0n 20n 70n)
Vcin 7 0 PULSE (0 5 0n 0n 0n 15n 70n)
.tran 1n 100n
.control
run
display
plot V(1) V(2) V(7)
plot V(11) V(12)
.endc
.end
