* opamp subcircuit
.subckt opamp 1 2 4 5
R1 1 2 2MEG
R2 3 5 75
Ea 4 3 1 2 2E+5
.ends opamp
