*opamp differentiator
.include opamp.cir
Xdiv1 2 0 0 3 opamp
Rf 2 3 2k
C1 1 2 1u
Vin 1 0 sin(0 1 1k)
.tran 10u 1m
.control
run
display
plot V(1) V(3)
.endc
.end
