*opamp differentiator practical
.include opamp.cir
Xdiv1 3 4 0 5 opamp
Rf 3 5 20k
r1 2 3 10k
r2 4 0 6.67k
C1 1 2 1n
Vin 1 0 PULSE (0 5 0n 0n 0n 45n 70n)
.tran 10n 100n
.control
run
display
plot V(1) V(5)
.endc
.end
